module fsm_mealy(clk, reset, en, xin, zout);
input clk, reset, en, xin;
output zout;

reg zout;


endmodule

