module  ha(a, b, sum, cout);
input a, b;
output sum, cout;




endmodule
