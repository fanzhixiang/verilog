module matrix_mul_test;

parameter CYCLE = 20;

parameter a = 7;
parameter b = 13;
parameter c = 5;




endmodule
