module STI(clk ,reset, load, pi_data,  pi_msb, pi_low,
           so_data, so_valid );

input       clk, reset;
input       load, pi_msb, pi_low; 
input   [15:0]  pi_data;

output      so_data, so_valid;





endmodule




