module fa(a, b, ci, sum, cout);
input  a, b, ci;
output sum, cout;




endmodule
