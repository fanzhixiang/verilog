module alu(alu_out, accum, data, opcode, zero, clk, reset);
input clk, reset;
input [7:0] accum, data;
input [2:0] opcode;
output [7:0] alu_out;
output zero;






endmodule
